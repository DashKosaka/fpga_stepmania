// DE2_115_SOPC.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		input  wire        Terasic_IrDA_0_conduit_end_export,                                                 //             Terasic_IrDA_0_conduit_end.export
		output wire        altpll_audio_locked_conduit_export,                                                //            altpll_audio_locked_conduit.export
		output wire        altpll_audio_phasedone_conduit_export,                                             //         altpll_audio_phasedone_conduit.export
		output wire        altpll_c1_clk,                                                                     //                              altpll_c1.clk
		output wire        altpll_c2_clk,                                                                     //                              altpll_c2.clk
		output wire        altpll_c3_clk,                                                                     //                              altpll_c3.clk
		output wire        altpll_c4_clk,                                                                     //                              altpll_c4.clk
		output wire        altpll_locked_conduit_export,                                                      //                  altpll_locked_conduit.export
		output wire        altpll_phasedone_conduit_export,                                                   //               altpll_phasedone_conduit.export
		output wire        audio_conduit_end_XCK,                                                             //                      audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                                                          //                                       .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                                                          //                                       .ADCLRC
		output wire        audio_conduit_end_DACDAT,                                                          //                                       .DACDAT
		input  wire        audio_conduit_end_DACLRC,                                                          //                                       .DACLRC
		input  wire        audio_conduit_end_BCLK,                                                            //                                       .BCLK
		input  wire        clk_50_clk_in_clk,                                                                 //                          clk_50_clk_in.clk
		input  wire        clk_50_clk_in_reset_reset_n,                                                       //                    clk_50_clk_in_reset.reset_n
		output wire        eep_i2c_scl_external_connection_export,                                            //        eep_i2c_scl_external_connection.export
		inout  wire        eep_i2c_sda_external_connection_export,                                            //        eep_i2c_sda_external_connection.export
		output wire        i2c_scl_external_connection_export,                                                //            i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,                                                //            i2c_sda_external_connection.export
		input  wire [3:0]  key_external_connection_export,                                                    //                key_external_connection.export
		output wire        lcd_external_RS,                                                                   //                           lcd_external.RS
		output wire        lcd_external_RW,                                                                   //                                       .RW
		inout  wire [7:0]  lcd_external_data,                                                                 //                                       .data
		output wire        lcd_external_E,                                                                    //                                       .E
		output wire [8:0]  ledg_external_connection_export,                                                   //               ledg_external_connection.export
		output wire [17:0] ledr_external_connection_export,                                                   //               ledr_external_connection.export
		input  wire        rs232_external_connection_rxd,                                                     //              rs232_external_connection.rxd
		output wire        rs232_external_connection_txd,                                                     //                                       .txd
		input  wire        rs232_external_connection_cts_n,                                                   //                                       .cts_n
		output wire        rs232_external_connection_rts_n,                                                   //                                       .rts_n
		output wire        sd_clk_external_connection_export,                                                 //             sd_clk_external_connection.export
		inout  wire        sd_cmd_external_connection_export,                                                 //             sd_cmd_external_connection.export
		inout  wire [3:0]  sd_dat_external_connection_export,                                                 //             sd_dat_external_connection.export
		input  wire        sd_wp_n_external_connection_export,                                                //            sd_wp_n_external_connection.export
		output wire [63:0] seg7_conduit_end_export,                                                           //                       seg7_conduit_end.export
		input  wire        sma_in_external_connection_export,                                                 //             sma_in_external_connection.export
		output wire        sma_out_external_connection_export,                                                //            sma_out_external_connection.export
		input  wire [17:0] sw_external_connection_export,                                                     //                 sw_external_connection.export
		output wire [22:0] tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_address_out,      // tri_state_bridge_flash_bridge_0_export.av_tri_s1_cfi_flash_0_tcm_address_out
		output wire [0:0]  tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_write_n_out,      //                                       .av_tri_s1_cfi_flash_0_tcm_write_n_out
		output wire [0:0]  tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out, //                                       .av_tri_s1_cfi_flash_0_tcm_chipselect_n_out
		output wire [0:0]  tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_read_n_out,       //                                       .av_tri_s1_cfi_flash_0_tcm_read_n_out
		inout  wire [7:0]  tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_data_out          //                                       .av_tri_s1_cfi_flash_0_tcm_data_out
	);

	wire         altpll_c0_clk;                                                                    // altpll:c0 -> [av_tri_s1_cfi_flash_0:clk_clk, clock_crossing_io:m0_clk, clock_crossing_io:s0_clk, cpu:clk, eep_i2c_scl:clk, eep_i2c_sda:clk, i2c_scl:clk, i2c_sda:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, key:clk, lcd:clk, ledg:clk, ledr:clk, mm_interconnect_0:altpll_c0_clk, mm_interconnect_1:altpll_c0_clk, onchip_memory2:clk, rs232:clk, rst_controller_002:clk, sd_clk:clk, sd_cmd:clk, sd_dat:clk, sd_wp_n:clk, seg7:s_clk, sma_in:clk, sma_out:clk, sw:clk, sysid:clock, timer:clk, tri_state_bridge_flash_bridge_0:clk, tristate_conduit_pin_sharer_0:clk_clk]
	wire         altpll_audio_c0_clk;                                                              // altpll_audio:c0 -> [audio:avs_s1_clk, mm_interconnect_0:altpll_audio_c0_clk, rst_controller_001:clk]
	wire   [7:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_in;          // tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_data_in -> tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_data_in
	wire         tristate_conduit_pin_sharer_0_tcm_request;                                        // tristate_conduit_pin_sharer_0:request -> tri_state_bridge_flash_bridge_0:request
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_write_n_out_out;      // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_write_n_out -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_write_n_out
	wire  [22:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_address_out_out;      // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_address_out -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_address_out
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_read_n_out_out;       // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_read_n_out -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_read_n_out
	wire         tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_outen;       // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_data_outen -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_data_outen
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out_out; // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_chipselect_n_out -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out
	wire         tristate_conduit_pin_sharer_0_tcm_grant;                                          // tri_state_bridge_flash_bridge_0:grant -> tristate_conduit_pin_sharer_0:grant
	wire   [7:0] tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_out;         // tristate_conduit_pin_sharer_0:av_tri_s1_cfi_flash_0_tcm_data_out -> tri_state_bridge_flash_bridge_0:tcs_av_tri_s1_cfi_flash_0_tcm_data_out
	wire         av_tri_s1_cfi_flash_0_tcm_data_outen;                                             // av_tri_s1_cfi_flash_0:tcm_data_outen -> tristate_conduit_pin_sharer_0:tcs0_data_outen
	wire         av_tri_s1_cfi_flash_0_tcm_request;                                                // av_tri_s1_cfi_flash_0:tcm_request -> tristate_conduit_pin_sharer_0:tcs0_request
	wire         av_tri_s1_cfi_flash_0_tcm_write_n_out;                                            // av_tri_s1_cfi_flash_0:tcm_write_n_out -> tristate_conduit_pin_sharer_0:tcs0_write_n_out
	wire         av_tri_s1_cfi_flash_0_tcm_read_n_out;                                             // av_tri_s1_cfi_flash_0:tcm_read_n_out -> tristate_conduit_pin_sharer_0:tcs0_read_n_out
	wire         av_tri_s1_cfi_flash_0_tcm_grant;                                                  // tristate_conduit_pin_sharer_0:tcs0_grant -> av_tri_s1_cfi_flash_0:tcm_grant
	wire         av_tri_s1_cfi_flash_0_tcm_chipselect_n_out;                                       // av_tri_s1_cfi_flash_0:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_0:tcs0_chipselect_n_out
	wire  [22:0] av_tri_s1_cfi_flash_0_tcm_address_out;                                            // av_tri_s1_cfi_flash_0:tcm_address_out -> tristate_conduit_pin_sharer_0:tcs0_address_out
	wire   [7:0] av_tri_s1_cfi_flash_0_tcm_data_out;                                               // av_tri_s1_cfi_flash_0:tcm_data_out -> tristate_conduit_pin_sharer_0:tcs0_data_out
	wire   [7:0] av_tri_s1_cfi_flash_0_tcm_data_in;                                                // tristate_conduit_pin_sharer_0:tcs0_data_in -> av_tri_s1_cfi_flash_0:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                                         // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                      // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                      // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                                          // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                       // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                             // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                                    // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                            // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                        // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                  // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                               // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                                                   // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                      // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                             // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_readdata;                                    // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_audio_avalon_slave_address;                                     // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire         mm_interconnect_0_audio_avalon_slave_read;                                        // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire         mm_interconnect_0_audio_avalon_slave_write;                                       // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_writedata;                                   // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire         mm_interconnect_0_terasic_irda_0_avalon_slave_chipselect;                         // mm_interconnect_0:Terasic_IrDA_0_avalon_slave_chipselect -> Terasic_IrDA_0:s_cs_n
	wire  [31:0] mm_interconnect_0_terasic_irda_0_avalon_slave_readdata;                           // Terasic_IrDA_0:s_readdata -> mm_interconnect_0:Terasic_IrDA_0_avalon_slave_readdata
	wire         mm_interconnect_0_terasic_irda_0_avalon_slave_read;                               // mm_interconnect_0:Terasic_IrDA_0_avalon_slave_read -> Terasic_IrDA_0:s_read
	wire         mm_interconnect_0_terasic_irda_0_avalon_slave_write;                              // mm_interconnect_0:Terasic_IrDA_0_avalon_slave_write -> Terasic_IrDA_0:s_write
	wire  [31:0] mm_interconnect_0_terasic_irda_0_avalon_slave_writedata;                          // mm_interconnect_0:Terasic_IrDA_0_avalon_slave_writedata -> Terasic_IrDA_0:s_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                   // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                    // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                       // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                 // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                      // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                  // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                                      // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                                       // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                                          // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                                         // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;                                     // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_readdata;                                // altpll_audio:readdata -> mm_interconnect_0:altpll_audio_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_audio_pll_slave_address;                                 // mm_interconnect_0:altpll_audio_pll_slave_address -> altpll_audio:address
	wire         mm_interconnect_0_altpll_audio_pll_slave_read;                                    // mm_interconnect_0:altpll_audio_pll_slave_read -> altpll_audio:read
	wire         mm_interconnect_0_altpll_audio_pll_slave_write;                                   // mm_interconnect_0:altpll_audio_pll_slave_write -> altpll_audio:write
	wire  [31:0] mm_interconnect_0_altpll_audio_pll_slave_writedata;                               // mm_interconnect_0:altpll_audio_pll_slave_writedata -> altpll_audio:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                                  // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                               // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                               // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire   [8:0] mm_interconnect_0_clock_crossing_io_s0_address;                                   // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                                      // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                                // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                             // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                                     // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                                 // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                                // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                                   // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                                     // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;                                      // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                                   // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                                        // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                                    // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                                        // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire  [31:0] mm_interconnect_0_sma_in_s1_readdata;                                             // sma_in:readdata -> mm_interconnect_0:sma_in_s1_readdata
	wire   [1:0] mm_interconnect_0_sma_in_s1_address;                                              // mm_interconnect_0:sma_in_s1_address -> sma_in:address
	wire         mm_interconnect_0_sma_out_s1_chipselect;                                          // mm_interconnect_0:sma_out_s1_chipselect -> sma_out:chipselect
	wire  [31:0] mm_interconnect_0_sma_out_s1_readdata;                                            // sma_out:readdata -> mm_interconnect_0:sma_out_s1_readdata
	wire   [1:0] mm_interconnect_0_sma_out_s1_address;                                             // mm_interconnect_0:sma_out_s1_address -> sma_out:address
	wire         mm_interconnect_0_sma_out_s1_write;                                               // mm_interconnect_0:sma_out_s1_write -> sma_out:write_n
	wire  [31:0] mm_interconnect_0_sma_out_s1_writedata;                                           // mm_interconnect_0:sma_out_s1_writedata -> sma_out:writedata
	wire   [7:0] mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdata;                             // av_tri_s1_cfi_flash_0:uas_readdata -> mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_readdata
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_waitrequest;                          // av_tri_s1_cfi_flash_0:uas_waitrequest -> mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_waitrequest
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_debugaccess;                          // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_debugaccess -> av_tri_s1_cfi_flash_0:uas_debugaccess
	wire  [22:0] mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_address;                              // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_address -> av_tri_s1_cfi_flash_0:uas_address
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_read;                                 // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_read -> av_tri_s1_cfi_flash_0:uas_read
	wire   [0:0] mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_byteenable;                           // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_byteenable -> av_tri_s1_cfi_flash_0:uas_byteenable
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdatavalid;                        // av_tri_s1_cfi_flash_0:uas_readdatavalid -> mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_readdatavalid
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_lock;                                 // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_lock -> av_tri_s1_cfi_flash_0:uas_lock
	wire         mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_write;                                // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_write -> av_tri_s1_cfi_flash_0:uas_write
	wire   [7:0] mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_writedata;                            // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_writedata -> av_tri_s1_cfi_flash_0:uas_writedata
	wire   [0:0] mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_burstcount;                           // mm_interconnect_0:av_tri_s1_cfi_flash_0_uas_burstcount -> av_tri_s1_cfi_flash_0:uas_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                                 // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                                                    // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                                 // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [8:0] clock_crossing_io_m0_address;                                                     // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                                        // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                                                  // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                               // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                                                   // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                                       // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                                                  // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_readdata;                                     // seg7:s_readdata -> mm_interconnect_1:seg7_avalon_slave_readdata
	wire   [2:0] mm_interconnect_1_seg7_avalon_slave_address;                                      // mm_interconnect_1:seg7_avalon_slave_address -> seg7:s_address
	wire         mm_interconnect_1_seg7_avalon_slave_read;                                         // mm_interconnect_1:seg7_avalon_slave_read -> seg7:s_read
	wire         mm_interconnect_1_seg7_avalon_slave_write;                                        // mm_interconnect_1:seg7_avalon_slave_write -> seg7:s_write
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_writedata;                                    // mm_interconnect_1:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                                   // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                                    // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;                                     // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;                                      // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_read;                                         // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;                                // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_1_lcd_control_slave_write;                                        // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;                                    // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire         mm_interconnect_1_timer_s1_chipselect;                                            // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                              // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                               // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                                                 // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                             // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_1_key_s1_chipselect;                                              // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                                // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                                 // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                                                   // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                               // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                                               // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                                 // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                                  // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                                                    // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                                // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_1_ledg_s1_chipselect;                                             // mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_1_ledg_s1_readdata;                                               // ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	wire   [1:0] mm_interconnect_1_ledg_s1_address;                                                // mm_interconnect_1:ledg_s1_address -> ledg:address
	wire         mm_interconnect_1_ledg_s1_write;                                                  // mm_interconnect_1:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_1_ledg_s1_writedata;                                              // mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_1_ledr_s1_chipselect;                                             // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                                               // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                                                // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_write;                                                  // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                                              // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_1_rs232_s1_chipselect;                                            // mm_interconnect_1:rs232_s1_chipselect -> rs232:chipselect
	wire  [15:0] mm_interconnect_1_rs232_s1_readdata;                                              // rs232:readdata -> mm_interconnect_1:rs232_s1_readdata
	wire   [2:0] mm_interconnect_1_rs232_s1_address;                                               // mm_interconnect_1:rs232_s1_address -> rs232:address
	wire         mm_interconnect_1_rs232_s1_read;                                                  // mm_interconnect_1:rs232_s1_read -> rs232:read_n
	wire         mm_interconnect_1_rs232_s1_begintransfer;                                         // mm_interconnect_1:rs232_s1_begintransfer -> rs232:begintransfer
	wire         mm_interconnect_1_rs232_s1_write;                                                 // mm_interconnect_1:rs232_s1_write -> rs232:write_n
	wire  [15:0] mm_interconnect_1_rs232_s1_writedata;                                             // mm_interconnect_1:rs232_s1_writedata -> rs232:writedata
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                                          // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                                            // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                                             // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_write;                                               // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                                           // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                                          // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                                            // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                                             // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_write;                                               // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                                           // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire         mm_interconnect_1_eep_i2c_scl_s1_chipselect;                                      // mm_interconnect_1:eep_i2c_scl_s1_chipselect -> eep_i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_eep_i2c_scl_s1_readdata;                                        // eep_i2c_scl:readdata -> mm_interconnect_1:eep_i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_eep_i2c_scl_s1_address;                                         // mm_interconnect_1:eep_i2c_scl_s1_address -> eep_i2c_scl:address
	wire         mm_interconnect_1_eep_i2c_scl_s1_write;                                           // mm_interconnect_1:eep_i2c_scl_s1_write -> eep_i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_eep_i2c_scl_s1_writedata;                                       // mm_interconnect_1:eep_i2c_scl_s1_writedata -> eep_i2c_scl:writedata
	wire         mm_interconnect_1_eep_i2c_sda_s1_chipselect;                                      // mm_interconnect_1:eep_i2c_sda_s1_chipselect -> eep_i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_eep_i2c_sda_s1_readdata;                                        // eep_i2c_sda:readdata -> mm_interconnect_1:eep_i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_eep_i2c_sda_s1_address;                                         // mm_interconnect_1:eep_i2c_sda_s1_address -> eep_i2c_sda:address
	wire         mm_interconnect_1_eep_i2c_sda_s1_write;                                           // mm_interconnect_1:eep_i2c_sda_s1_write -> eep_i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_eep_i2c_sda_s1_writedata;                                       // mm_interconnect_1:eep_i2c_sda_s1_writedata -> eep_i2c_sda:writedata
	wire         mm_interconnect_1_sd_clk_s1_chipselect;                                           // mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	wire  [31:0] mm_interconnect_1_sd_clk_s1_readdata;                                             // sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_clk_s1_address;                                              // mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	wire         mm_interconnect_1_sd_clk_s1_write;                                                // mm_interconnect_1:sd_clk_s1_write -> sd_clk:write_n
	wire  [31:0] mm_interconnect_1_sd_clk_s1_writedata;                                            // mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	wire         mm_interconnect_1_sd_cmd_s1_chipselect;                                           // mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_readdata;                                             // sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_cmd_s1_address;                                              // mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	wire         mm_interconnect_1_sd_cmd_s1_write;                                                // mm_interconnect_1:sd_cmd_s1_write -> sd_cmd:write_n
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_writedata;                                            // mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	wire         mm_interconnect_1_sd_dat_s1_chipselect;                                           // mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	wire  [31:0] mm_interconnect_1_sd_dat_s1_readdata;                                             // sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_dat_s1_address;                                              // mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	wire         mm_interconnect_1_sd_dat_s1_write;                                                // mm_interconnect_1:sd_dat_s1_write -> sd_dat:write_n
	wire  [31:0] mm_interconnect_1_sd_dat_s1_writedata;                                            // mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	wire  [31:0] mm_interconnect_1_sd_wp_n_s1_readdata;                                            // sd_wp_n:readdata -> mm_interconnect_1:sd_wp_n_s1_readdata
	wire   [1:0] mm_interconnect_1_sd_wp_n_s1_address;                                             // mm_interconnect_1:sd_wp_n_s1_address -> sd_wp_n:address
	wire         irq_mapper_receiver1_irq;                                                         // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                         // key:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                         // sw:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                         // rs232:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                         // jtag_uart:av_irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_irq_irq;                                                                      // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver0_irq;                                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                    // Terasic_IrDA_0:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [Terasic_IrDA_0:reset_n, altpll:reset, altpll_audio:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                               // rst_controller_001:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_clock_sink_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                               // rst_controller_002:reset_out -> [av_tri_s1_cfi_flash_0:reset_reset, clock_crossing_io:m0_reset, clock_crossing_io:s0_reset, cpu:reset_n, eep_i2c_scl:reset_n, eep_i2c_sda:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, key:reset_n, lcd:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rs232:reset_n, rst_translator:in_reset, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, sd_wp_n:reset_n, seg7:s_reset, sma_in:reset_n, sma_out:reset_n, sw:reset_n, sysid:reset_n, timer:reset_n, tri_state_bridge_flash_bridge_0:reset, tristate_conduit_pin_sharer_0:reset_reset]
	wire         rst_controller_002_reset_out_reset_req;                                           // rst_controller_002:reset_req -> [cpu:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]

	TERASIC_IRM terasic_irda_0 (
		.s_read      (mm_interconnect_0_terasic_irda_0_avalon_slave_read),        //     avalon_slave.read
		.s_cs_n      (~mm_interconnect_0_terasic_irda_0_avalon_slave_chipselect), //                 .chipselect_n
		.s_readdata  (mm_interconnect_0_terasic_irda_0_avalon_slave_readdata),    //                 .readdata
		.s_write     (mm_interconnect_0_terasic_irda_0_avalon_slave_write),       //                 .write
		.s_writedata (mm_interconnect_0_terasic_irda_0_avalon_slave_writedata),   //                 .writedata
		.clk         (clk_50_clk_in_clk),                                         //       clock_sink.clk
		.reset_n     (~rst_controller_reset_out_reset),                           // clock_sink_reset.reset_n
		.ir          (Terasic_IrDA_0_conduit_end_export),                         //      conduit_end.export
		.irq         (irq_synchronizer_receiver_irq)                              // interrupt_sender.irq
	);

	DE2_115_SOPC_altpll altpll (
		.clk       (clk_50_clk_in_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                //                    c0.clk
		.c1        (altpll_c1_clk),                                //                    c1.clk
		.c2        (altpll_c2_clk),                                //                    c2.clk
		.c3        (altpll_c3_clk),                                //                    c3.clk
		.c4        (altpll_c4_clk),                                //                    c4.clk
		.areset    (),                                             //        areset_conduit.export
		.locked    (altpll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	DE2_115_SOPC_altpll_audio altpll_audio (
		.clk       (clk_50_clk_in_clk),                                  //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                     // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_audio_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_audio_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_audio_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_audio_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_audio_pll_slave_writedata), //                      .writedata
		.c0        (altpll_audio_c0_clk),                                //                    c0.clk
		.locked    (altpll_audio_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_audio_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	AUDIO_IF audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (altpll_audio_c0_clk),                            //       clock_sink.clk
		.avs_s1_reset         (rst_controller_001_reset_out_reset),             // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	DE2_115_SOPC_av_tri_s1_cfi_flash_0 #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) av_tri_s1_cfi_flash_0 (
		.clk_clk              (altpll_c0_clk),                                             //   clk.clk
		.reset_reset          (rst_controller_002_reset_out_reset),                        // reset.reset
		.uas_address          (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (av_tri_s1_cfi_flash_0_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (av_tri_s1_cfi_flash_0_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (av_tri_s1_cfi_flash_0_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (av_tri_s1_cfi_flash_0_tcm_request),                         //      .request
		.tcm_grant            (av_tri_s1_cfi_flash_0_tcm_grant),                           //      .grant
		.tcm_address_out      (av_tri_s1_cfi_flash_0_tcm_address_out),                     //      .address_out
		.tcm_data_out         (av_tri_s1_cfi_flash_0_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (av_tri_s1_cfi_flash_0_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (av_tri_s1_cfi_flash_0_tcm_data_in)                          //      .data_in
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_c0_clk),                                        //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (altpll_c0_clk),                                        //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                 (altpll_c0_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DE2_115_SOPC_eep_i2c_scl eep_i2c_scl (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_eep_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_eep_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_eep_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_eep_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_eep_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (eep_i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_eep_i2c_sda eep_i2c_sda (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_eep_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_eep_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_eep_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_eep_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_eep_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (eep_i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_eep_i2c_scl i2c_scl (
		.clk        (altpll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_eep_i2c_sda i2c_sda (
		.clk        (altpll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver5_irq)                                   //               irq.irq
	);

	DE2_115_SOPC_key key (
		.clk        (altpll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	DE2_115_SOPC_lcd lcd (
		.reset_n       (~rst_controller_002_reset_out_reset),               //         reset.reset_n
		.clk           (altpll_c0_clk),                                     //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_external_RS),                                   //      external.export
		.LCD_RW        (lcd_external_RW),                                   //              .export
		.LCD_data      (lcd_external_data),                                 //              .export
		.LCD_E         (lcd_external_E)                                     //              .export
	);

	DE2_115_SOPC_ledg ledg (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_ledr ledr (
		.clk        (altpll_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_onchip_memory2 onchip_memory2 (
		.clk        (altpll_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)          //       .reset_req
	);

	DE2_115_SOPC_rs232 rs232 (
		.clk           (altpll_c0_clk),                            //                 clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address       (mm_interconnect_1_rs232_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_rs232_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_rs232_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_rs232_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_rs232_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_rs232_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_rs232_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (rs232_external_connection_rxd),            // external_connection.export
		.txd           (rs232_external_connection_txd),            //                    .export
		.cts_n         (rs232_external_connection_cts_n),          //                    .export
		.rts_n         (rs232_external_connection_rts_n),          //                    .export
		.irq           (irq_mapper_receiver4_irq)                  //                 irq.irq
	);

	DE2_115_SOPC_eep_i2c_scl sd_clk (
		.clk        (altpll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_eep_i2c_sda sd_cmd (
		.clk        (altpll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sd_dat sd_dat (
		.clk        (altpll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sd_wp_n sd_wp_n (
		.clk      (altpll_c0_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_1_sd_wp_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sd_wp_n_s1_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)     // external_connection.export
	);

	SEG7_IF #(
		.SEG7_NUM       (8),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_1_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_1_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_1_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_1_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_1_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                       //      conduit_end.export
		.s_clk       (altpll_c0_clk),                                 //       clock_sink.clk
		.s_reset     (rst_controller_002_reset_out_reset)             // clock_sink_reset.reset
	);

	DE2_115_SOPC_sd_wp_n sma_in (
		.clk      (altpll_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sma_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sma_in_s1_readdata), //                    .readdata
		.in_port  (sma_in_external_connection_export)     // external_connection.export
	);

	DE2_115_SOPC_eep_i2c_scl sma_out (
		.clk        (altpll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_sma_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sma_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sma_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sma_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sma_out_s1_readdata),   //                    .readdata
		.out_port   (sma_out_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sw sw (
		.clk        (altpll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_mapper_receiver3_irq)             //                 irq.irq
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_timer timer (
		.clk        (altpll_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	DE2_115_SOPC_tri_state_bridge_flash_bridge_0 tri_state_bridge_flash_bridge_0 (
		.clk                                            (altpll_c0_clk),                                                                     //   clk.clk
		.reset                                          (rst_controller_002_reset_out_reset),                                                // reset.reset
		.request                                        (tristate_conduit_pin_sharer_0_tcm_request),                                         //   tcs.request
		.grant                                          (tristate_conduit_pin_sharer_0_tcm_grant),                                           //      .grant
		.tcs_av_tri_s1_cfi_flash_0_tcm_address_out      (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_address_out_out),       //      .av_tri_s1_cfi_flash_0_tcm_address_out_out
		.tcs_av_tri_s1_cfi_flash_0_tcm_write_n_out      (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_write_n_out_out),       //      .av_tri_s1_cfi_flash_0_tcm_write_n_out_out
		.tcs_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out_out),  //      .av_tri_s1_cfi_flash_0_tcm_chipselect_n_out_out
		.tcs_av_tri_s1_cfi_flash_0_tcm_read_n_out       (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_read_n_out_out),        //      .av_tri_s1_cfi_flash_0_tcm_read_n_out_out
		.tcs_av_tri_s1_cfi_flash_0_tcm_data_out         (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_out),          //      .av_tri_s1_cfi_flash_0_tcm_data_out_out
		.tcs_av_tri_s1_cfi_flash_0_tcm_data_outen       (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_outen),        //      .av_tri_s1_cfi_flash_0_tcm_data_out_outen
		.tcs_av_tri_s1_cfi_flash_0_tcm_data_in          (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_in),           //      .av_tri_s1_cfi_flash_0_tcm_data_out_in
		.av_tri_s1_cfi_flash_0_tcm_address_out          (tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_address_out),      //   out.av_tri_s1_cfi_flash_0_tcm_address_out
		.av_tri_s1_cfi_flash_0_tcm_write_n_out          (tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_write_n_out),      //      .av_tri_s1_cfi_flash_0_tcm_write_n_out
		.av_tri_s1_cfi_flash_0_tcm_chipselect_n_out     (tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out), //      .av_tri_s1_cfi_flash_0_tcm_chipselect_n_out
		.av_tri_s1_cfi_flash_0_tcm_read_n_out           (tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_read_n_out),       //      .av_tri_s1_cfi_flash_0_tcm_read_n_out
		.av_tri_s1_cfi_flash_0_tcm_data_out             (tri_state_bridge_flash_bridge_0_export_av_tri_s1_cfi_flash_0_tcm_data_out)          //      .av_tri_s1_cfi_flash_0_tcm_data_out
	);

	DE2_115_SOPC_tristate_conduit_pin_sharer_0 tristate_conduit_pin_sharer_0 (
		.clk_clk                                    (altpll_c0_clk),                                                                    //   clk.clk
		.reset_reset                                (rst_controller_002_reset_out_reset),                                               // reset.reset
		.request                                    (tristate_conduit_pin_sharer_0_tcm_request),                                        //   tcm.request
		.grant                                      (tristate_conduit_pin_sharer_0_tcm_grant),                                          //      .grant
		.av_tri_s1_cfi_flash_0_tcm_address_out      (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_address_out_out),      //      .av_tri_s1_cfi_flash_0_tcm_address_out_out
		.av_tri_s1_cfi_flash_0_tcm_read_n_out       (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_read_n_out_out),       //      .av_tri_s1_cfi_flash_0_tcm_read_n_out_out
		.av_tri_s1_cfi_flash_0_tcm_write_n_out      (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_write_n_out_out),      //      .av_tri_s1_cfi_flash_0_tcm_write_n_out_out
		.av_tri_s1_cfi_flash_0_tcm_data_out         (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_out),         //      .av_tri_s1_cfi_flash_0_tcm_data_out_out
		.av_tri_s1_cfi_flash_0_tcm_data_in          (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_in),          //      .av_tri_s1_cfi_flash_0_tcm_data_out_in
		.av_tri_s1_cfi_flash_0_tcm_data_outen       (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_data_out_outen),       //      .av_tri_s1_cfi_flash_0_tcm_data_out_outen
		.av_tri_s1_cfi_flash_0_tcm_chipselect_n_out (tristate_conduit_pin_sharer_0_tcm_av_tri_s1_cfi_flash_0_tcm_chipselect_n_out_out), //      .av_tri_s1_cfi_flash_0_tcm_chipselect_n_out_out
		.tcs0_request                               (av_tri_s1_cfi_flash_0_tcm_request),                                                //  tcs0.request
		.tcs0_grant                                 (av_tri_s1_cfi_flash_0_tcm_grant),                                                  //      .grant
		.tcs0_address_out                           (av_tri_s1_cfi_flash_0_tcm_address_out),                                            //      .address_out
		.tcs0_read_n_out                            (av_tri_s1_cfi_flash_0_tcm_read_n_out),                                             //      .read_n_out
		.tcs0_write_n_out                           (av_tri_s1_cfi_flash_0_tcm_write_n_out),                                            //      .write_n_out
		.tcs0_data_out                              (av_tri_s1_cfi_flash_0_tcm_data_out),                                               //      .data_out
		.tcs0_data_in                               (av_tri_s1_cfi_flash_0_tcm_data_in),                                                //      .data_in
		.tcs0_data_outen                            (av_tri_s1_cfi_flash_0_tcm_data_outen),                                             //      .data_outen
		.tcs0_chipselect_n_out                      (av_tri_s1_cfi_flash_0_tcm_chipselect_n_out)                                        //      .chipselect_n_out
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                             //                                          altpll_c0.clk
		.altpll_audio_c0_clk                                      (altpll_audio_c0_clk),                                       //                                    altpll_audio_c0.clk
		.clk_50_clk_clk                                           (clk_50_clk_in_clk),                                         //                                         clk_50_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.audio_clock_sink_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                        //       audio_clock_sink_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                    (rst_controller_002_reset_out_reset),                        //                    cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                  (cpu_data_master_address),                                   //                                    cpu_data_master.address
		.cpu_data_master_waitrequest                              (cpu_data_master_waitrequest),                               //                                                   .waitrequest
		.cpu_data_master_byteenable                               (cpu_data_master_byteenable),                                //                                                   .byteenable
		.cpu_data_master_read                                     (cpu_data_master_read),                                      //                                                   .read
		.cpu_data_master_readdata                                 (cpu_data_master_readdata),                                  //                                                   .readdata
		.cpu_data_master_readdatavalid                            (cpu_data_master_readdatavalid),                             //                                                   .readdatavalid
		.cpu_data_master_write                                    (cpu_data_master_write),                                     //                                                   .write
		.cpu_data_master_writedata                                (cpu_data_master_writedata),                                 //                                                   .writedata
		.cpu_data_master_debugaccess                              (cpu_data_master_debugaccess),                               //                                                   .debugaccess
		.cpu_instruction_master_address                           (cpu_instruction_master_address),                            //                             cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                       (cpu_instruction_master_waitrequest),                        //                                                   .waitrequest
		.cpu_instruction_master_read                              (cpu_instruction_master_read),                               //                                                   .read
		.cpu_instruction_master_readdata                          (cpu_instruction_master_readdata),                           //                                                   .readdata
		.cpu_instruction_master_readdatavalid                     (cpu_instruction_master_readdatavalid),                      //                                                   .readdatavalid
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                  //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                   //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),               //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),              //                                                   .writedata
		.altpll_audio_pll_slave_address                           (mm_interconnect_0_altpll_audio_pll_slave_address),          //                             altpll_audio_pll_slave.address
		.altpll_audio_pll_slave_write                             (mm_interconnect_0_altpll_audio_pll_slave_write),            //                                                   .write
		.altpll_audio_pll_slave_read                              (mm_interconnect_0_altpll_audio_pll_slave_read),             //                                                   .read
		.altpll_audio_pll_slave_readdata                          (mm_interconnect_0_altpll_audio_pll_slave_readdata),         //                                                   .readdata
		.altpll_audio_pll_slave_writedata                         (mm_interconnect_0_altpll_audio_pll_slave_writedata),        //                                                   .writedata
		.audio_avalon_slave_address                               (mm_interconnect_0_audio_avalon_slave_address),              //                                 audio_avalon_slave.address
		.audio_avalon_slave_write                                 (mm_interconnect_0_audio_avalon_slave_write),                //                                                   .write
		.audio_avalon_slave_read                                  (mm_interconnect_0_audio_avalon_slave_read),                 //                                                   .read
		.audio_avalon_slave_readdata                              (mm_interconnect_0_audio_avalon_slave_readdata),             //                                                   .readdata
		.audio_avalon_slave_writedata                             (mm_interconnect_0_audio_avalon_slave_writedata),            //                                                   .writedata
		.av_tri_s1_cfi_flash_0_uas_address                        (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_address),       //                          av_tri_s1_cfi_flash_0_uas.address
		.av_tri_s1_cfi_flash_0_uas_write                          (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_write),         //                                                   .write
		.av_tri_s1_cfi_flash_0_uas_read                           (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_read),          //                                                   .read
		.av_tri_s1_cfi_flash_0_uas_readdata                       (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdata),      //                                                   .readdata
		.av_tri_s1_cfi_flash_0_uas_writedata                      (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_writedata),     //                                                   .writedata
		.av_tri_s1_cfi_flash_0_uas_burstcount                     (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_burstcount),    //                                                   .burstcount
		.av_tri_s1_cfi_flash_0_uas_byteenable                     (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_byteenable),    //                                                   .byteenable
		.av_tri_s1_cfi_flash_0_uas_readdatavalid                  (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_readdatavalid), //                                                   .readdatavalid
		.av_tri_s1_cfi_flash_0_uas_waitrequest                    (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_waitrequest),   //                                                   .waitrequest
		.av_tri_s1_cfi_flash_0_uas_lock                           (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_lock),          //                                                   .lock
		.av_tri_s1_cfi_flash_0_uas_debugaccess                    (mm_interconnect_0_av_tri_s1_cfi_flash_0_uas_debugaccess),   //                                                   .debugaccess
		.clock_crossing_io_s0_address                             (mm_interconnect_0_clock_crossing_io_s0_address),            //                               clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                               (mm_interconnect_0_clock_crossing_io_s0_write),              //                                                   .write
		.clock_crossing_io_s0_read                                (mm_interconnect_0_clock_crossing_io_s0_read),               //                                                   .read
		.clock_crossing_io_s0_readdata                            (mm_interconnect_0_clock_crossing_io_s0_readdata),           //                                                   .readdata
		.clock_crossing_io_s0_writedata                           (mm_interconnect_0_clock_crossing_io_s0_writedata),          //                                                   .writedata
		.clock_crossing_io_s0_burstcount                          (mm_interconnect_0_clock_crossing_io_s0_burstcount),         //                                                   .burstcount
		.clock_crossing_io_s0_byteenable                          (mm_interconnect_0_clock_crossing_io_s0_byteenable),         //                                                   .byteenable
		.clock_crossing_io_s0_readdatavalid                       (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),      //                                                   .readdatavalid
		.clock_crossing_io_s0_waitrequest                         (mm_interconnect_0_clock_crossing_io_s0_waitrequest),        //                                                   .waitrequest
		.clock_crossing_io_s0_debugaccess                         (mm_interconnect_0_clock_crossing_io_s0_debugaccess),        //                                                   .debugaccess
		.cpu_debug_mem_slave_address                              (mm_interconnect_0_cpu_debug_mem_slave_address),             //                                cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                                   .write
		.cpu_debug_mem_slave_read                                 (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                                   .read
		.cpu_debug_mem_slave_readdata                             (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                                   .readdata
		.cpu_debug_mem_slave_writedata                            (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                                   .writedata
		.cpu_debug_mem_slave_byteenable                           (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                                   .byteenable
		.cpu_debug_mem_slave_waitrequest                          (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                                   .waitrequest
		.cpu_debug_mem_slave_debugaccess                          (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                                   .debugaccess
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                   .chipselect
		.onchip_memory2_s1_address                                (mm_interconnect_0_onchip_memory2_s1_address),               //                                  onchip_memory2_s1.address
		.onchip_memory2_s1_write                                  (mm_interconnect_0_onchip_memory2_s1_write),                 //                                                   .write
		.onchip_memory2_s1_readdata                               (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                                   .readdata
		.onchip_memory2_s1_writedata                              (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                                   .writedata
		.onchip_memory2_s1_byteenable                             (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                                   .byteenable
		.onchip_memory2_s1_chipselect                             (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                                   .chipselect
		.onchip_memory2_s1_clken                                  (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                                   .clken
		.sma_in_s1_address                                        (mm_interconnect_0_sma_in_s1_address),                       //                                          sma_in_s1.address
		.sma_in_s1_readdata                                       (mm_interconnect_0_sma_in_s1_readdata),                      //                                                   .readdata
		.sma_out_s1_address                                       (mm_interconnect_0_sma_out_s1_address),                      //                                         sma_out_s1.address
		.sma_out_s1_write                                         (mm_interconnect_0_sma_out_s1_write),                        //                                                   .write
		.sma_out_s1_readdata                                      (mm_interconnect_0_sma_out_s1_readdata),                     //                                                   .readdata
		.sma_out_s1_writedata                                     (mm_interconnect_0_sma_out_s1_writedata),                    //                                                   .writedata
		.sma_out_s1_chipselect                                    (mm_interconnect_0_sma_out_s1_chipselect),                   //                                                   .chipselect
		.Terasic_IrDA_0_avalon_slave_write                        (mm_interconnect_0_terasic_irda_0_avalon_slave_write),       //                        Terasic_IrDA_0_avalon_slave.write
		.Terasic_IrDA_0_avalon_slave_read                         (mm_interconnect_0_terasic_irda_0_avalon_slave_read),        //                                                   .read
		.Terasic_IrDA_0_avalon_slave_readdata                     (mm_interconnect_0_terasic_irda_0_avalon_slave_readdata),    //                                                   .readdata
		.Terasic_IrDA_0_avalon_slave_writedata                    (mm_interconnect_0_terasic_irda_0_avalon_slave_writedata),   //                                                   .writedata
		.Terasic_IrDA_0_avalon_slave_chipselect                   (mm_interconnect_0_terasic_irda_0_avalon_slave_chipselect)   //                                                   .chipselect
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.altpll_c0_clk                                          (altpll_c0_clk),                                     //                                        altpll_c0.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                      //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                  //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                   //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                   //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                         //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                     //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                        //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                    //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                  //                                                 .debugaccess
		.eep_i2c_scl_s1_address                                 (mm_interconnect_1_eep_i2c_scl_s1_address),          //                                   eep_i2c_scl_s1.address
		.eep_i2c_scl_s1_write                                   (mm_interconnect_1_eep_i2c_scl_s1_write),            //                                                 .write
		.eep_i2c_scl_s1_readdata                                (mm_interconnect_1_eep_i2c_scl_s1_readdata),         //                                                 .readdata
		.eep_i2c_scl_s1_writedata                               (mm_interconnect_1_eep_i2c_scl_s1_writedata),        //                                                 .writedata
		.eep_i2c_scl_s1_chipselect                              (mm_interconnect_1_eep_i2c_scl_s1_chipselect),       //                                                 .chipselect
		.eep_i2c_sda_s1_address                                 (mm_interconnect_1_eep_i2c_sda_s1_address),          //                                   eep_i2c_sda_s1.address
		.eep_i2c_sda_s1_write                                   (mm_interconnect_1_eep_i2c_sda_s1_write),            //                                                 .write
		.eep_i2c_sda_s1_readdata                                (mm_interconnect_1_eep_i2c_sda_s1_readdata),         //                                                 .readdata
		.eep_i2c_sda_s1_writedata                               (mm_interconnect_1_eep_i2c_sda_s1_writedata),        //                                                 .writedata
		.eep_i2c_sda_s1_chipselect                              (mm_interconnect_1_eep_i2c_sda_s1_chipselect),       //                                                 .chipselect
		.i2c_scl_s1_address                                     (mm_interconnect_1_i2c_scl_s1_address),              //                                       i2c_scl_s1.address
		.i2c_scl_s1_write                                       (mm_interconnect_1_i2c_scl_s1_write),                //                                                 .write
		.i2c_scl_s1_readdata                                    (mm_interconnect_1_i2c_scl_s1_readdata),             //                                                 .readdata
		.i2c_scl_s1_writedata                                   (mm_interconnect_1_i2c_scl_s1_writedata),            //                                                 .writedata
		.i2c_scl_s1_chipselect                                  (mm_interconnect_1_i2c_scl_s1_chipselect),           //                                                 .chipselect
		.i2c_sda_s1_address                                     (mm_interconnect_1_i2c_sda_s1_address),              //                                       i2c_sda_s1.address
		.i2c_sda_s1_write                                       (mm_interconnect_1_i2c_sda_s1_write),                //                                                 .write
		.i2c_sda_s1_readdata                                    (mm_interconnect_1_i2c_sda_s1_readdata),             //                                                 .readdata
		.i2c_sda_s1_writedata                                   (mm_interconnect_1_i2c_sda_s1_writedata),            //                                                 .writedata
		.i2c_sda_s1_chipselect                                  (mm_interconnect_1_i2c_sda_s1_chipselect),           //                                                 .chipselect
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),                  //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                    //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),                 //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),                //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),               //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),       //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),         //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),          //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),      //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),     //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer), //                                                 .begintransfer
		.ledg_s1_address                                        (mm_interconnect_1_ledg_s1_address),                 //                                          ledg_s1.address
		.ledg_s1_write                                          (mm_interconnect_1_ledg_s1_write),                   //                                                 .write
		.ledg_s1_readdata                                       (mm_interconnect_1_ledg_s1_readdata),                //                                                 .readdata
		.ledg_s1_writedata                                      (mm_interconnect_1_ledg_s1_writedata),               //                                                 .writedata
		.ledg_s1_chipselect                                     (mm_interconnect_1_ledg_s1_chipselect),              //                                                 .chipselect
		.ledr_s1_address                                        (mm_interconnect_1_ledr_s1_address),                 //                                          ledr_s1.address
		.ledr_s1_write                                          (mm_interconnect_1_ledr_s1_write),                   //                                                 .write
		.ledr_s1_readdata                                       (mm_interconnect_1_ledr_s1_readdata),                //                                                 .readdata
		.ledr_s1_writedata                                      (mm_interconnect_1_ledr_s1_writedata),               //                                                 .writedata
		.ledr_s1_chipselect                                     (mm_interconnect_1_ledr_s1_chipselect),              //                                                 .chipselect
		.rs232_s1_address                                       (mm_interconnect_1_rs232_s1_address),                //                                         rs232_s1.address
		.rs232_s1_write                                         (mm_interconnect_1_rs232_s1_write),                  //                                                 .write
		.rs232_s1_read                                          (mm_interconnect_1_rs232_s1_read),                   //                                                 .read
		.rs232_s1_readdata                                      (mm_interconnect_1_rs232_s1_readdata),               //                                                 .readdata
		.rs232_s1_writedata                                     (mm_interconnect_1_rs232_s1_writedata),              //                                                 .writedata
		.rs232_s1_begintransfer                                 (mm_interconnect_1_rs232_s1_begintransfer),          //                                                 .begintransfer
		.rs232_s1_chipselect                                    (mm_interconnect_1_rs232_s1_chipselect),             //                                                 .chipselect
		.sd_clk_s1_address                                      (mm_interconnect_1_sd_clk_s1_address),               //                                        sd_clk_s1.address
		.sd_clk_s1_write                                        (mm_interconnect_1_sd_clk_s1_write),                 //                                                 .write
		.sd_clk_s1_readdata                                     (mm_interconnect_1_sd_clk_s1_readdata),              //                                                 .readdata
		.sd_clk_s1_writedata                                    (mm_interconnect_1_sd_clk_s1_writedata),             //                                                 .writedata
		.sd_clk_s1_chipselect                                   (mm_interconnect_1_sd_clk_s1_chipselect),            //                                                 .chipselect
		.sd_cmd_s1_address                                      (mm_interconnect_1_sd_cmd_s1_address),               //                                        sd_cmd_s1.address
		.sd_cmd_s1_write                                        (mm_interconnect_1_sd_cmd_s1_write),                 //                                                 .write
		.sd_cmd_s1_readdata                                     (mm_interconnect_1_sd_cmd_s1_readdata),              //                                                 .readdata
		.sd_cmd_s1_writedata                                    (mm_interconnect_1_sd_cmd_s1_writedata),             //                                                 .writedata
		.sd_cmd_s1_chipselect                                   (mm_interconnect_1_sd_cmd_s1_chipselect),            //                                                 .chipselect
		.sd_dat_s1_address                                      (mm_interconnect_1_sd_dat_s1_address),               //                                        sd_dat_s1.address
		.sd_dat_s1_write                                        (mm_interconnect_1_sd_dat_s1_write),                 //                                                 .write
		.sd_dat_s1_readdata                                     (mm_interconnect_1_sd_dat_s1_readdata),              //                                                 .readdata
		.sd_dat_s1_writedata                                    (mm_interconnect_1_sd_dat_s1_writedata),             //                                                 .writedata
		.sd_dat_s1_chipselect                                   (mm_interconnect_1_sd_dat_s1_chipselect),            //                                                 .chipselect
		.sd_wp_n_s1_address                                     (mm_interconnect_1_sd_wp_n_s1_address),              //                                       sd_wp_n_s1.address
		.sd_wp_n_s1_readdata                                    (mm_interconnect_1_sd_wp_n_s1_readdata),             //                                                 .readdata
		.seg7_avalon_slave_address                              (mm_interconnect_1_seg7_avalon_slave_address),       //                                seg7_avalon_slave.address
		.seg7_avalon_slave_write                                (mm_interconnect_1_seg7_avalon_slave_write),         //                                                 .write
		.seg7_avalon_slave_read                                 (mm_interconnect_1_seg7_avalon_slave_read),          //                                                 .read
		.seg7_avalon_slave_readdata                             (mm_interconnect_1_seg7_avalon_slave_readdata),      //                                                 .readdata
		.seg7_avalon_slave_writedata                            (mm_interconnect_1_seg7_avalon_slave_writedata),     //                                                 .writedata
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                   //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                     //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),                  //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),                 //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),                //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),     //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata),    //                                                 .readdata
		.timer_s1_address                                       (mm_interconnect_1_timer_s1_address),                //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_1_timer_s1_write),                  //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_1_timer_s1_readdata),               //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_1_timer_s1_writedata),              //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_1_timer_s1_chipselect)              //                                                 .chipselect
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_50_clk_in_clk),                  //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_50_clk_in_reset_reset_n),   // reset_in0.reset
		.clk            (clk_50_clk_in_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_50_clk_in_reset_reset_n),       // reset_in0.reset
		.clk            (altpll_audio_c0_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~clk_50_clk_in_reset_reset_n),           // reset_in0.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
