module step_chart(
	input logic Clk, reset, frame_clk,
	output logic [3:0] display_signal
);


logic [3:0] step_chart[100]='{4'b1111, 
										   4'b0000,
										   4'b1010,
										   4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0101,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1010,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1001,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0110,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0101,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1010,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1001,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0110,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0101,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1010,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1001,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0110,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0101,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1010,
											4'b0000,
											4'b0000,
											4'b0101,
                                 4'b0000,
                                 4'b0000,
											4'b0000,
											4'b0000,
											4'b0000,
											4'b1010,
											4'b0000
											};
											
											
											
											
											
											
											
//bit [3:0] step_chart[2:0];// = [4'b1010, 4'b0000];
/*
parameter [399:0] step_chart = { {4'b0101}, 
										   {4'b0000},
										   {4'b1010},
										   {4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0101},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1010},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1001},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0110},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0101},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1010},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1001},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0110},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0101},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1010},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1001},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0110},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0101},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b0000},
											{4'b1010},
											{4'b0000}
											};
*/
										  
										  
//parameter [3:0] step_chart [2] = 4'b0000;
//step_chart [1][3:0] = 4'b0000;
/*
parameter [3:0] step_chart[1:100] ={4'b1010,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0101,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1010,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1001,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0110,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0101,											
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1010,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1001,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0110,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0101,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1010,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1001,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0110,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0101,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1010,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b1001,
												4'b0000,
												4'b0000,
												4'b0000,
												4'b0000};
 */                                      
//step_chart[1] = 42;                  
                                       
logic frame_clk_delayed;
logic frame_clk_rising_edge;

logic [8:0] current, next;

always_ff @ (posedge Clk)
begin
    frame_clk_delayed <= frame_clk;
end
assign frame_clk_rising_edge = (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);

always_ff @ (posedge Clk)
begin
    if(reset)
    begin
		step_chart <='{4'b1111, 
							4'b0000,
							4'b1010,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0101,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1010,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1001,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0110,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0101,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1010,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1001,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0110,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0101,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1010,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1001,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0110,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0101,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1010,
							4'b0000,
							4'b0000,
							4'b0101,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b0000,
							4'b1010,
							4'b0000
							};
    end
    else if(frame_clk_rising_edge)
    begin
		//current <= next;
		display_signal <= step_chart[1];
//		step_chart <= 4'b1010;
		for(int i=1;i<99;i++)
		begin
			step_chart[i-1] <= step_chart[i];
		end
	 end
end
/*
always_comb
begin

	next = current + 9'h4;
	if(current + 9'h4 > 9'h399)
	begin
		next = 9'b0;
	end

end
*/
endmodule